`default_nettype none
`timescale 1ns/1ps

/*
this testbench just instantiates the module and makes some convenient wires
that can be driven / tested by the cocotb test.py
*/

// testbench is controlled by test.py
module tb (
    // system
    input   clk,
    input   rst_n,
    input   ena,
    // spi
    input   spi_sck,
    input   spi_sce,
    input   spi_sin,
    output  spi_sout,
    // adc spi
    output  adc_sck,
    output  adc_sce,
    input   adc_sin,
    output  adc_sout
);

    // this part dumps the trace to a vcd file that can be viewed with GTKWave
    initial begin
        $dumpfile ("tb.vcd");
        $dumpvars (0, tb);
        `ifndef VERILATOR
            #1;
        `endif
    end

    wire [7:0] ui_in = { 4'b0, adc_sin, spi_sin, spi_sce, spi_sck };
    wire [7:0] uo_out;
    wire [7:0] uio_in = 8'b0;
    wire [7:0] uio_out;
    wire [7:0] uio_oe;
    assign { adc_sout, adc_sce, adc_sck, spi_sout } = uo_out[3:0];

    tt_um_thermocouple tt_um_thermocouple (
    // include power ports for the Gate Level test
    `ifdef GL_TEST
        .VPWR( 1'b1),
        .VGND( 1'b0),
    `endif
        .ui_in      (ui_in),    // Dedicated inputs
        .uo_out     (uo_out),   // Dedicated outputs
        .uio_in     (uio_in),   // IOs: Input path
        .uio_out    (uio_out),  // IOs: Output path
        .uio_oe     (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
        .ena        (ena),      // enable - goes high when design is selected
        .clk        (clk),      // clock
        .rst_n      (rst_n)     // not reset
    );

endmodule
